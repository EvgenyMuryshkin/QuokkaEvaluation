`default_nettype none

module CombinationalROMModule_TopLevel (
	input  [7: 0] ReadAddress1,
	input  [7: 0] ReadAddress2,
	output [7: 0] Value1,
	output [7: 0] Value2
    );

reg [7:0] MemoryBlock [0 : 255];
initial
begin
	MemoryBlock[0] = 8'b00011111;
	MemoryBlock[1] = 8'b00101011;
	MemoryBlock[2] = 8'b11010011;
	MemoryBlock[3] = 8'b11101101;
	MemoryBlock[4] = 8'b11010010;
	MemoryBlock[5] = 8'b11100101;
	MemoryBlock[6] = 8'b01101011;
	MemoryBlock[7] = 8'b01110010;
	MemoryBlock[8] = 8'b10111111;
	MemoryBlock[9] = 8'b11101101;
	MemoryBlock[10] = 8'b01011111;
	MemoryBlock[11] = 8'b01100010;
	MemoryBlock[12] = 8'b10010000;
	MemoryBlock[13] = 8'b10011010;
	MemoryBlock[14] = 8'b11101110;
	MemoryBlock[15] = 8'b00010000;
	MemoryBlock[16] = 8'b11000000;
	MemoryBlock[17] = 8'b10111011;
	MemoryBlock[18] = 8'b01001010;
	MemoryBlock[19] = 8'b01101000;
	MemoryBlock[20] = 8'b00101111;
	MemoryBlock[21] = 8'b10100110;
	MemoryBlock[22] = 8'b01000111;
	MemoryBlock[23] = 8'b01010000;
	MemoryBlock[24] = 8'b00000000;
	MemoryBlock[25] = 8'b00100100;
	MemoryBlock[26] = 8'b10011001;
	MemoryBlock[27] = 8'b01010100;
	MemoryBlock[28] = 8'b01011101;
	MemoryBlock[29] = 8'b10100110;
	MemoryBlock[30] = 8'b10110011;
	MemoryBlock[31] = 8'b01110011;
	MemoryBlock[32] = 8'b01011111;
	MemoryBlock[33] = 8'b01111011;
	MemoryBlock[34] = 8'b11000011;
	MemoryBlock[35] = 8'b00110000;
	MemoryBlock[36] = 8'b01101011;
	MemoryBlock[37] = 8'b11001111;
	MemoryBlock[38] = 8'b11011110;
	MemoryBlock[39] = 8'b01000000;
	MemoryBlock[40] = 8'b11101100;
	MemoryBlock[41] = 8'b01101100;
	MemoryBlock[42] = 8'b00101011;
	MemoryBlock[43] = 8'b00000001;
	MemoryBlock[44] = 8'b01010111;
	MemoryBlock[45] = 8'b10010011;
	MemoryBlock[46] = 8'b11111000;
	MemoryBlock[47] = 8'b01000110;
	MemoryBlock[48] = 8'b00100010;
	MemoryBlock[49] = 8'b01000001;
	MemoryBlock[50] = 8'b10110100;
	MemoryBlock[51] = 8'b01100100;
	MemoryBlock[52] = 8'b11011010;
	MemoryBlock[53] = 8'b10010110;
	MemoryBlock[54] = 8'b01000111;
	MemoryBlock[55] = 8'b01111000;
	MemoryBlock[56] = 8'b11100011;
	MemoryBlock[57] = 8'b10000010;
	MemoryBlock[58] = 8'b11101100;
	MemoryBlock[59] = 8'b10101101;
	MemoryBlock[60] = 8'b01001100;
	MemoryBlock[61] = 8'b00010111;
	MemoryBlock[62] = 8'b00010100;
	MemoryBlock[63] = 8'b00011000;
	MemoryBlock[64] = 8'b00111010;
	MemoryBlock[65] = 8'b11101011;
	MemoryBlock[66] = 8'b00000011;
	MemoryBlock[67] = 8'b00010101;
	MemoryBlock[68] = 8'b11010110;
	MemoryBlock[69] = 8'b10111101;
	MemoryBlock[70] = 8'b10100101;
	MemoryBlock[71] = 8'b11110000;
	MemoryBlock[72] = 8'b11011100;
	MemoryBlock[73] = 8'b00001010;
	MemoryBlock[74] = 8'b01111011;
	MemoryBlock[75] = 8'b11000010;
	MemoryBlock[76] = 8'b01111010;
	MemoryBlock[77] = 8'b01000110;
	MemoryBlock[78] = 8'b11111001;
	MemoryBlock[79] = 8'b01101100;
	MemoryBlock[80] = 8'b00101011;
	MemoryBlock[81] = 8'b01010010;
	MemoryBlock[82] = 8'b00110001;
	MemoryBlock[83] = 8'b00011100;
	MemoryBlock[84] = 8'b11110010;
	MemoryBlock[85] = 8'b01001110;
	MemoryBlock[86] = 8'b10011000;
	MemoryBlock[87] = 8'b11001001;
	MemoryBlock[88] = 8'b00110011;
	MemoryBlock[89] = 8'b01001010;
	MemoryBlock[90] = 8'b01001100;
	MemoryBlock[91] = 8'b11101001;
	MemoryBlock[92] = 8'b11100010;
	MemoryBlock[93] = 8'b00110001;
	MemoryBlock[94] = 8'b11110011;
	MemoryBlock[95] = 8'b11010101;
	MemoryBlock[96] = 8'b01011000;
	MemoryBlock[97] = 8'b00010010;
	MemoryBlock[98] = 8'b11000110;
	MemoryBlock[99] = 8'b01101011;
	MemoryBlock[100] = 8'b10010000;
	MemoryBlock[101] = 8'b11100011;
	MemoryBlock[102] = 8'b01110000;
	MemoryBlock[103] = 8'b01100100;
	MemoryBlock[104] = 8'b10011100;
	MemoryBlock[105] = 8'b11000011;
	MemoryBlock[106] = 8'b10000111;
	MemoryBlock[107] = 8'b11010000;
	MemoryBlock[108] = 8'b00011010;
	MemoryBlock[109] = 8'b10000101;
	MemoryBlock[110] = 8'b11111110;
	MemoryBlock[111] = 8'b10011101;
	MemoryBlock[112] = 8'b10001000;
	MemoryBlock[113] = 8'b01111111;
	MemoryBlock[114] = 8'b10000001;
	MemoryBlock[115] = 8'b11111001;
	MemoryBlock[116] = 8'b11100101;
	MemoryBlock[117] = 8'b11111000;
	MemoryBlock[118] = 8'b00100110;
	MemoryBlock[119] = 8'b11101011;
	MemoryBlock[120] = 8'b01010011;
	MemoryBlock[121] = 8'b00111001;
	MemoryBlock[122] = 8'b11100001;
	MemoryBlock[123] = 8'b10001011;
	MemoryBlock[124] = 8'b01110001;
	MemoryBlock[125] = 8'b10111011;
	MemoryBlock[126] = 8'b00001110;
	MemoryBlock[127] = 8'b10101011;
	MemoryBlock[128] = 8'b00010110;
	MemoryBlock[129] = 8'b10100110;
	MemoryBlock[130] = 8'b01101010;
	MemoryBlock[131] = 8'b01100111;
	MemoryBlock[132] = 8'b01111111;
	MemoryBlock[133] = 8'b10001110;
	MemoryBlock[134] = 8'b11011100;
	MemoryBlock[135] = 8'b01000111;
	MemoryBlock[136] = 8'b11100010;
	MemoryBlock[137] = 8'b11001101;
	MemoryBlock[138] = 8'b10000000;
	MemoryBlock[139] = 8'b00101110;
	MemoryBlock[140] = 8'b11000110;
	MemoryBlock[141] = 8'b11000111;
	MemoryBlock[142] = 8'b10101110;
	MemoryBlock[143] = 8'b10101110;
	MemoryBlock[144] = 8'b01001100;
	MemoryBlock[145] = 8'b10101110;
	MemoryBlock[146] = 8'b01100000;
	MemoryBlock[147] = 8'b01100011;
	MemoryBlock[148] = 8'b10101111;
	MemoryBlock[149] = 8'b11111001;
	MemoryBlock[150] = 8'b11101111;
	MemoryBlock[151] = 8'b01011111;
	MemoryBlock[152] = 8'b11101100;
	MemoryBlock[153] = 8'b11011011;
	MemoryBlock[154] = 8'b00011000;
	MemoryBlock[155] = 8'b01010110;
	MemoryBlock[156] = 8'b00000010;
	MemoryBlock[157] = 8'b11100100;
	MemoryBlock[158] = 8'b11110011;
	MemoryBlock[159] = 8'b11100000;
	MemoryBlock[160] = 8'b10110101;
	MemoryBlock[161] = 8'b11011011;
	MemoryBlock[162] = 8'b10111010;
	MemoryBlock[163] = 8'b01110011;
	MemoryBlock[164] = 8'b00011010;
	MemoryBlock[165] = 8'b10010110;
	MemoryBlock[166] = 8'b00011110;
	MemoryBlock[167] = 8'b11111010;
	MemoryBlock[168] = 8'b10100011;
	MemoryBlock[169] = 8'b00111001;
	MemoryBlock[170] = 8'b00010111;
	MemoryBlock[171] = 8'b00011000;
	MemoryBlock[172] = 8'b01111000;
	MemoryBlock[173] = 8'b11111000;
	MemoryBlock[174] = 8'b00100100;
	MemoryBlock[175] = 8'b10001011;
	MemoryBlock[176] = 8'b10001010;
	MemoryBlock[177] = 8'b00110011;
	MemoryBlock[178] = 8'b00111111;
	MemoryBlock[179] = 8'b11000010;
	MemoryBlock[180] = 8'b01011010;
	MemoryBlock[181] = 8'b10101011;
	MemoryBlock[182] = 8'b11111100;
	MemoryBlock[183] = 8'b00011100;
	MemoryBlock[184] = 8'b10110110;
	MemoryBlock[185] = 8'b00001010;
	MemoryBlock[186] = 8'b01111011;
	MemoryBlock[187] = 8'b10100100;
	MemoryBlock[188] = 8'b01110110;
	MemoryBlock[189] = 8'b10000101;
	MemoryBlock[190] = 8'b01000101;
	MemoryBlock[191] = 8'b11111110;
	MemoryBlock[192] = 8'b11011001;
	MemoryBlock[193] = 8'b10011111;
	MemoryBlock[194] = 8'b01111001;
	MemoryBlock[195] = 8'b11101011;
	MemoryBlock[196] = 8'b00001100;
	MemoryBlock[197] = 8'b00111010;
	MemoryBlock[198] = 8'b10010011;
	MemoryBlock[199] = 8'b10110101;
	MemoryBlock[200] = 8'b10010000;
	MemoryBlock[201] = 8'b01100110;
	MemoryBlock[202] = 8'b10111111;
	MemoryBlock[203] = 8'b01110101;
	MemoryBlock[204] = 8'b11100010;
	MemoryBlock[205] = 8'b11010111;
	MemoryBlock[206] = 8'b11100111;
	MemoryBlock[207] = 8'b11110100;
	MemoryBlock[208] = 8'b10110110;
	MemoryBlock[209] = 8'b10001100;
	MemoryBlock[210] = 8'b11001011;
	MemoryBlock[211] = 8'b11001111;
	MemoryBlock[212] = 8'b10100101;
	MemoryBlock[213] = 8'b00110001;
	MemoryBlock[214] = 8'b10000101;
	MemoryBlock[215] = 8'b00001010;
	MemoryBlock[216] = 8'b11011111;
	MemoryBlock[217] = 8'b10011110;
	MemoryBlock[218] = 8'b10111100;
	MemoryBlock[219] = 8'b00001111;
	MemoryBlock[220] = 8'b00011011;
	MemoryBlock[221] = 8'b01111001;
	MemoryBlock[222] = 8'b10000011;
	MemoryBlock[223] = 8'b00011110;
	MemoryBlock[224] = 8'b11110100;
	MemoryBlock[225] = 8'b00011001;
	MemoryBlock[226] = 8'b00111110;
	MemoryBlock[227] = 8'b11011000;
	MemoryBlock[228] = 8'b01111110;
	MemoryBlock[229] = 8'b00111001;
	MemoryBlock[230] = 8'b01111111;
	MemoryBlock[231] = 8'b01010000;
	MemoryBlock[232] = 8'b10011111;
	MemoryBlock[233] = 8'b10001001;
	MemoryBlock[234] = 8'b00110001;
	MemoryBlock[235] = 8'b11110100;
	MemoryBlock[236] = 8'b11101011;
	MemoryBlock[237] = 8'b10000111;
	MemoryBlock[238] = 8'b00111001;
	MemoryBlock[239] = 8'b11011111;
	MemoryBlock[240] = 8'b00100010;
	MemoryBlock[241] = 8'b10000111;
	MemoryBlock[242] = 8'b11101110;
	MemoryBlock[243] = 8'b11101010;
	MemoryBlock[244] = 8'b10111001;
	MemoryBlock[245] = 8'b01110101;
	MemoryBlock[246] = 8'b01011000;
	MemoryBlock[247] = 8'b10101000;
	MemoryBlock[248] = 8'b00011001;
	MemoryBlock[249] = 8'b01101111;
	MemoryBlock[250] = 8'b00001011;
	MemoryBlock[251] = 8'b01101110;
	MemoryBlock[252] = 8'b01111101;
	MemoryBlock[253] = 8'b10000011;
	MemoryBlock[254] = 8'b10011010;
	MemoryBlock[255] = 8'b00010110;
end

assign Value1 = MemoryBlock[ReadAddress1];
assign Value2 = MemoryBlock[ReadAddress2];

endmodule
